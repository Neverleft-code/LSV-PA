module top(o, a, b, c);
output o;
input a, b, c;
//wire t_0, t_1, t_2;
and g1(o, a, b, c);
endmodule
